// haze-cpu: decoder_5to32.sv
// (c) 2025 Connor J. Link. All rights reserved.

module decoder_5to32
(
    input  logic [4:0]  i_S,
    output logic [31:0] o_Q
);

    always_comb begin
        unique case (i_S)
            5'b00000: o_Q = 32'b00000000000000000000000000000001;
            5'b00001: o_Q = 32'b00000000000000000000000000000010;
            5'b00010: o_Q = 32'b00000000000000000000000000000100;
            5'b00011: o_Q = 32'b00000000000000000000000000001000;
            5'b00100: o_Q = 32'b00000000000000000000000000010000;
            5'b00101: o_Q = 32'b00000000000000000000000000100000;
            5'b00110: o_Q = 32'b00000000000000000000000001000000;
            5'b00111: o_Q = 32'b00000000000000000000000010000000;
            5'b01000: o_Q = 32'b00000000000000000000000100000000;
            5'b01001: o_Q = 32'b00000000000000000000001000000000;
            5'b01010: o_Q = 32'b00000000000000000000010000000000;
            5'b01011: o_Q = 32'b00000000000000000000100000000000;
            5'b01100: o_Q = 32'b00000000000000000001000000000000;
            5'b01101: o_Q = 32'b00000000000000000010000000000000;
            5'b01110: o_Q = 32'b00000000000000000100000000000000;
            5'b01111: o_Q = 32'b00000000000000001000000000000000;
            5'b10000: o_Q = 32'b00000000000000010000000000000000;
            5'b10001: o_Q = 32'b00000000000000100000000000000000;
            5'b10010: o_Q = 32'b00000000000001000000000000000000;
            5'b10011: o_Q = 32'b00000000000010000000000000000000;
            5'b10100: o_Q = 32'b00000000000100000000000000000000;
            5'b10101: o_Q = 32'b00000000001000000000000000000000;
            5'b10110: o_Q = 32'b00000000010000000000000000000000;
            5'b10111: o_Q = 32'b00000000100000000000000000000000;
            5'b11000: o_Q = 32'b00000001000000000000000000000000;
            5'b11001: o_Q = 32'b00000010000000000000000000000000;
            5'b11010: o_Q = 32'b00000100000000000000000000000000;
            5'b11011: o_Q = 32'b00001000000000000000000000000000;
            5'b11100: o_Q = 32'b00010000000000000000000000000000;
            5'b11101: o_Q = 32'b00100000000000000000000000000000;
            5'b11110: o_Q = 32'b01000000000000000000000000000000;
            5'b11111: o_Q = 32'b10000000000000000000000000000000;
            default:  o_Q = 32'b00000000000000000000000000000000; // fallback
        endcase
    end

endmodule