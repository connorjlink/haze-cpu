-- Horizon: register_IF.vhd
-- (c) 2026 Connor J. Link. All rights reserved.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.types.all;

entity register_IF is
    port(
        i_Clock    : in  std_logic;
        i_Reset    : in  std_logic;
        i_Stall    : in  std_logic;
        i_Flush    : in  std_logic;
        i_Signals  : in  IF_record_t;
        o_Signals  : out IF_record_t
    );
end register_IF;

architecture implementation of register_IF is
begin

    g_PipelineRegister: entity work.pipeline_register
        generic map(
            T   => IF_record_t,
            NOP => IF_NOP
        )
        port map(
            i_Clock   => i_Clock,
            i_Reset   => i_Reset,
            i_Stall   => i_Stall,
            i_Flush   => i_Flush,
            i_Signals => i_Signals,
            o_Signals => o_Signals
        );

end implementation;
